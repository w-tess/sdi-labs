library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb_butterfly is
end entity tb_butterfly;

architecture test of tb_butterfly is
	
begin
	
	
	
end architecture test;