library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity butterfly is
	port (
		
	);
end entity butterfly;

architecture behavioral of butterfly is
	
begin
	
	
	
end architecture behavioral;