library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fft_1616 is

end entity fft_1616;

architecture behavioral of fft_1616 is
	
begin
	
	
	
end architecture behavioral;